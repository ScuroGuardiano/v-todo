module utils

pub struct ApiError {
pub:
  error string
  status_code int
}
