module dto

pub struct TodoDtoDelete {
pub:
  id i64
}
